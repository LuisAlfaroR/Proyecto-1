
module AND( input wire ent1,ent2,output wire sal
    );

assign sal=ent1&ent2;

endmodule
